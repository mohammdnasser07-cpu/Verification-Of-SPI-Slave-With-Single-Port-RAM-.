package shared_pkg_slave;

endpackage