package shared_pkg;

endpackage